module top_module ( input x, input y, output z );
    xnor(z, x, y);
endmodule
